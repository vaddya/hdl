module lab2_4(a, res);

input [1:0] a;
output [5:0] res = a ** 3;

endmodule

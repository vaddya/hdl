module lab2_1(a, b, res);

input signed [3:0] a, b;
output signed [4:0] res = a + b;

endmodule

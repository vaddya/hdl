
module lab2_qsys (
	clk_clk,
	led_export,
	buttons_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	led_export;
	input		buttons_export;
	input		reset_reset_n;
endmodule

module lab2_2(a, b, res);

input signed [3:0] a, b;
output signed [6:0] res = a * b;

endmodule

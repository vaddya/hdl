module elab2_2(a, res);

input signed [3:0] a;
output signed [7:0] res = a * 9;

endmodule
